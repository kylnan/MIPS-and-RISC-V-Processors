`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/13/2021 12:44:35 PM
// Design Name: 
// Module Name: data_memory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module data_memory(
    input clk,
    input [31:0] mem_access_addr,
    input [31:0] mem_write_data,
    input mem_write_en,
    input mem_read_en,
    output [31:0] mem_read_data);
  
    integer i;  
    reg [31:0] ram [255:0];  // Don't change this name
    wire [7 : 0] ram_addr = mem_access_addr[9 : 2];  
    
    initial 
    begin 
       for(i=0;i<256;i=i+1)  
           ram[i] <= 32'd0;     
    end  
        
    always @(posedge clk) 
    begin  
       if (mem_write_en)  
           ram[ram_addr] <= mem_write_data;
       ram[0] = 32'd0 << 2;
       ram[1] = 32'd500;
       ram[2] = 32'd10;
       ram[3] = 32'd243;
       
       ram[9] = 32'd9 << 2;
       ram[10] = 32'd289;
       ram[11] = 32'd321;
    end  
      
    assign mem_read_data = (mem_read_en==1'b1) ? ram[ram_addr]: 32'd0;
            
endmodule
